/*module numberToDigits(input number, output digit0, output digit1, output digit2, output digit3);
	
	input [7:0] number;
	
	output [3:0] digit0;
	output [3:0] digit1;
	output [3:0] digit2;
	output [3:0] digit3;
	
	
	

endmodule*/
